`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:54:38 09/17/2021 
// Design Name: 
// Module Name:    practice2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module practice2;

	reg[3:0] start, result;
	initial;
	begin;
		start = 1;
		result = (start<<2);
	end
endmodule
