module practice (
    input a,
    output wire b
);

assign b = a + 1'sb0;

endmodule //practice

localparam 