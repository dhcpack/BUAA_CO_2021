`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   21:14:18 10/12/2021
// Design Name:   full_adder
// Module Name:   E:/ISE/learn/learn20211012/full_addwe_tb.v
// Project Name:  learn20211012
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: full_adder
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module full_addwe_tb;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	full_adder uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

