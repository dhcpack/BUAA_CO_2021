module practice (
    initial
    begin
      $display("hello world");
      $finish
      end
  );
endmodule //practice